package Skeleton_package;

//=============================================================================
// 			PARAMETERS		
//=============================================================================
	parameter NUM_MASTERS = 4;
	parameter NUM_SLAVES = 2;


//=============================================================================
// 			ADDRESS MAP		
//=============================================================================

	parameter USB_IFace_OFFSET 	= 35840;
	parameter USB_IFace_SIZE 	= 1024; 


	parameter TEST_RAM_OFFSET = 8192;
	parameter TEST_RAM_SIZE = 256;


endpackage 