package Skeleton_package;

//=============================================================================
// 			PARAMETERS		
//=============================================================================
	parameter NUM_MASTERS = 1;
	parameter NUM_SLAVES = 1;


//=============================================================================
// 			ADDRESS MAP		
//=============================================================================

	parameter TEST_RAM_OFFSET = 4096;
	parameter TEST_RAM_SIZE = 256;


endpackage 